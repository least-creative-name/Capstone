Example netlist
R1 N002 N001 100
C1 N002 0 100f
V1 N001 0 AC 1
.ac dec 20 1000 1e8
.backanno
.end
