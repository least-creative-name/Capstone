Example netlist
v1 1 0 dc 15
r1 1 0 2k
r2 1 2 1k
r3 2 0 1k
.op
.end
